
module memory_S(
    input              clk,
	input 			   rst_n,
    input     [7:0]    addr ,
    output reg[7:0]    mem_out
);

(* ramstyle = "M9K" *)    reg [7:0]	int_mem_i [255:0];  //S盒

    reg [3:0] a;
    reg [3:0] b;
    reg [7:0] ad;

    always @( * ) begin
       a=addr[7:4];
       b=addr[3:0];
       ad=(a<<4)+b;

    end
    
    always@(posedge clk or negedge rst_n )  begin
		if(!rst_n) begin
                    int_mem_i [8'h00] <=  8'h63 ;
                    int_mem_i [8'h01] <=  8'h7c ;
                    int_mem_i [8'h02] <=  8'h77 ;
                    int_mem_i [8'h03] <=  8'h7b ;
                    int_mem_i [8'h04] <=  8'hf2 ;
                    int_mem_i [8'h05] <=  8'h6b ;
                    int_mem_i [8'h06] <=  8'h6f ;
                    int_mem_i [8'h07] <=  8'hc5 ;
                    int_mem_i [8'h08] <=  8'h30 ;
                    int_mem_i [8'h09] <=  8'h01 ;
                    int_mem_i [8'h0a] <=  8'h67 ;
                    int_mem_i [8'h0b] <=  8'h2b ;
                    int_mem_i [8'h0c] <=  8'hfe ;
                    int_mem_i [8'h0d] <=  8'hd7 ;
                    int_mem_i [8'h0e] <=  8'hab ;
                    int_mem_i [8'h0f] <=  8'h76 ;
                    int_mem_i [8'h10] <=  8'hca ;
                    int_mem_i [8'h11] <=  8'h82 ;
                    int_mem_i [8'h12] <=  8'hc9 ;
                    int_mem_i [8'h13] <=  8'h7d ;
                    int_mem_i [8'h14] <=  8'hfa ;
                    int_mem_i [8'h15] <=  8'h59 ;
                    int_mem_i [8'h16] <=  8'h47 ;
                    int_mem_i [8'h17] <=  8'hf0 ;
                    int_mem_i [8'h18] <=  8'had ;
                    int_mem_i [8'h19] <=  8'hd4 ;
                    int_mem_i [8'h1a] <=  8'ha2 ;
                    int_mem_i [8'h1b] <=  8'haf ;
                    int_mem_i [8'h1c] <=  8'h9c ;
                    int_mem_i [8'h1d] <=  8'ha4 ;
                    int_mem_i [8'h1e] <=  8'h72 ;
                    int_mem_i [8'h1f] <=  8'hc0 ;
                    int_mem_i [8'h20] <=  8'hb7 ;
                    int_mem_i [8'h21] <=  8'hfd ;
                    int_mem_i [8'h22] <=  8'h93 ;
                    int_mem_i [8'h23] <=  8'h26 ;
                    int_mem_i [8'h24] <=  8'h36 ;
                    int_mem_i [8'h25] <=  8'h3f ;
                    int_mem_i [8'h26] <=  8'hf7 ;
                    int_mem_i [8'h27] <=  8'hcc ;
                    int_mem_i [8'h28] <=  8'h34 ;
                    int_mem_i [8'h29] <=  8'ha5 ;
                    int_mem_i [8'h2a] <=  8'he5 ;
                    int_mem_i [8'h2b] <=  8'hf1 ;
                    int_mem_i [8'h2c] <=  8'h71 ;
                    int_mem_i [8'h2d] <=  8'hd8 ;
                    int_mem_i [8'h2e] <=  8'h31 ;
                    int_mem_i [8'h2f] <=  8'h15 ;
                    int_mem_i [8'h30] <=  8'h04 ;
                    int_mem_i [8'h31] <=  8'hc7 ;
                    int_mem_i [8'h32] <=  8'h23 ;
                    int_mem_i [8'h33] <=  8'hc3 ;
                    int_mem_i [8'h34] <=  8'h18 ;
                    int_mem_i [8'h35] <=  8'h96 ;
                    int_mem_i [8'h36] <=  8'h05 ;
                    int_mem_i [8'h37] <=  8'h9a ;
                    int_mem_i [8'h38] <=  8'h07 ;
                    int_mem_i [8'h39] <=  8'h12 ;
                    int_mem_i [8'h3a] <=  8'h80 ;
                    int_mem_i [8'h3b] <=  8'he2 ;
                    int_mem_i [8'h3c] <=  8'heb ;
                    int_mem_i [8'h3d] <=  8'h27 ;
                    int_mem_i [8'h3e] <=  8'hb2 ;
                    int_mem_i [8'h3f] <=  8'h75 ;
                    int_mem_i [8'h40] <=  8'h09 ;
                    int_mem_i [8'h41] <=  8'h83 ;
                    int_mem_i [8'h42] <=  8'h2c ;
                    int_mem_i [8'h43] <=  8'h1a ;
                    int_mem_i [8'h44] <=  8'h1b ;
                    int_mem_i [8'h45] <=  8'h6e ;
                    int_mem_i [8'h46] <=  8'h5a ;
                    int_mem_i [8'h47] <=  8'ha0 ;
                    int_mem_i [8'h48] <=  8'h52 ;
                    int_mem_i [8'h49] <=  8'h3b ;
                    int_mem_i [8'h4a] <=  8'hd6 ;
                    int_mem_i [8'h4b] <=  8'hb3 ;
                    int_mem_i [8'h4c] <=  8'h29 ;
                    int_mem_i [8'h4d] <=  8'he3 ;
                    int_mem_i [8'h4e] <=  8'h2f ;
                    int_mem_i [8'h4f] <=  8'h84 ;
                    int_mem_i [8'h50] <=  8'h53 ;
                    int_mem_i [8'h51] <=  8'hd1 ;
                    int_mem_i [8'h52] <=  8'h00 ;
                    int_mem_i [8'h53] <=  8'hed ;
                    int_mem_i [8'h54] <=  8'h20 ;
                    int_mem_i [8'h55] <=  8'hfc ;
                    int_mem_i [8'h56] <=  8'hb1 ;
                    int_mem_i [8'h57] <=  8'h5b ;
                    int_mem_i [8'h58] <=  8'h6a ;
                    int_mem_i [8'h59] <=  8'hcb ;
                    int_mem_i [8'h5a] <=  8'hbe ;
                    int_mem_i [8'h5b] <=  8'h39 ;
                    int_mem_i [8'h5c] <=  8'h4a ;
                    int_mem_i [8'h5d] <=  8'h4c ;
                    int_mem_i [8'h5e] <=  8'h58 ;
                    int_mem_i [8'h5f] <=  8'hcf ;
                    int_mem_i [8'h60] <=  8'hd0 ;
                    int_mem_i [8'h61] <=  8'hef ;
                    int_mem_i [8'h62] <=  8'haa ;
                    int_mem_i [8'h63] <=  8'hfb ;
                    int_mem_i [8'h64] <=  8'h43 ;
                    int_mem_i [8'h65] <=  8'h4d ;
                    int_mem_i [8'h66] <=  8'h33 ;
                    int_mem_i [8'h67] <=  8'h85 ;
                    int_mem_i [8'h68] <=  8'h45 ;
                    int_mem_i [8'h69] <=  8'hf9 ;
                    int_mem_i [8'h6a] <=  8'h02 ;
                    int_mem_i [8'h6b] <=  8'h7f ;
                    int_mem_i [8'h6c] <=  8'h50 ;
                    int_mem_i [8'h6d] <=  8'h3c ;
                    int_mem_i [8'h6e] <=  8'h9f ;
                    int_mem_i [8'h6f] <=  8'ha8 ;
                    int_mem_i [8'h70] <=  8'h51 ;
                    int_mem_i [8'h71] <=  8'ha3 ;
                    int_mem_i [8'h72] <=  8'h40 ;
                    int_mem_i [8'h73] <=  8'h8f ;
                    int_mem_i [8'h74] <=  8'h92 ;
                    int_mem_i [8'h75] <=  8'h9d ;
                    int_mem_i [8'h76] <=  8'h38 ;
                    int_mem_i [8'h77] <=  8'hf5 ;
                    int_mem_i [8'h78] <=  8'hbc ;
                    int_mem_i [8'h79] <=  8'hb6 ;
                    int_mem_i [8'h7a] <=  8'hda ;
                    int_mem_i [8'h7b] <=  8'h21 ;
                    int_mem_i [8'h7c] <=  8'h10 ;
                    int_mem_i [8'h7d] <=  8'hff ;
                    int_mem_i [8'h7e] <=  8'hf3 ;
                    int_mem_i [8'h7f] <=  8'hd2 ;
                    int_mem_i [8'h80] <=  8'hcd ;
                    int_mem_i [8'h81] <=  8'h0c ;
                    int_mem_i [8'h82] <=  8'h13 ;
                    int_mem_i [8'h83] <=  8'hec ;
                    int_mem_i [8'h84] <=  8'h5f ;
                    int_mem_i [8'h85] <=  8'h97 ;
                    int_mem_i [8'h86] <=  8'h44 ;
                    int_mem_i [8'h87] <=  8'h17 ;
                    int_mem_i [8'h88] <=  8'hc4 ;
                    int_mem_i [8'h89] <=  8'ha7 ;
                    int_mem_i [8'h8a] <=  8'h7e ;
                    int_mem_i [8'h8b] <=  8'h3d ;
                    int_mem_i [8'h8c] <=  8'h64 ;
                    int_mem_i [8'h8d] <=  8'h5d ;
                    int_mem_i [8'h8e] <=  8'h19 ;
                    int_mem_i [8'h8f] <=  8'h73 ;
                    int_mem_i [8'h90] <=  8'h60 ;
                    int_mem_i [8'h91] <=  8'h81 ;
                    int_mem_i [8'h92] <=  8'h4f ;
                    int_mem_i [8'h93] <=  8'hdc ;
                    int_mem_i [8'h94] <=  8'h22 ;
                    int_mem_i [8'h95] <=  8'h2a ;
                    int_mem_i [8'h96] <=  8'h90 ;
                    int_mem_i [8'h97] <=  8'h88 ;
                    int_mem_i [8'h98] <=  8'h46 ;
                    int_mem_i [8'h99] <=  8'hee ;
                    int_mem_i [8'h9a] <=  8'hb8 ;
                    int_mem_i [8'h9b] <=  8'h14 ;
                    int_mem_i [8'h9c] <=  8'hde ;
                    int_mem_i [8'h9d] <=  8'h5e ;
                    int_mem_i [8'h9e] <=  8'h0b ;
                    int_mem_i [8'h9f] <=  8'hdb ;
                    int_mem_i [8'ha0] <=  8'he0 ;
                    int_mem_i [8'ha1] <=  8'h32 ;
                    int_mem_i [8'ha2] <=  8'h3a ;
                    int_mem_i [8'ha3] <=  8'h0a ;
                    int_mem_i [8'ha4] <=  8'h49 ;
                    int_mem_i [8'ha5] <=  8'h06 ;
                    int_mem_i [8'ha6] <=  8'h24 ;
                    int_mem_i [8'ha7] <=  8'h5c ;
                    int_mem_i [8'ha8] <=  8'hc2 ;
                    int_mem_i [8'ha9] <=  8'hd3 ;
                    int_mem_i [8'haa] <=  8'hac ;
                    int_mem_i [8'hab] <=  8'h62 ;
                    int_mem_i [8'hac] <=  8'h91 ;
                    int_mem_i [8'had] <=  8'h95 ;
                    int_mem_i [8'hae] <=  8'he4 ;
                    int_mem_i [8'haf] <=  8'h79 ;
                    int_mem_i [8'hb0] <=  8'he7 ;
                    int_mem_i [8'hb1] <=  8'hc8 ;
                    int_mem_i [8'hb2] <=  8'h37 ;
                    int_mem_i [8'hb3] <=  8'h6d ;
                    int_mem_i [8'hb4] <=  8'h8d ;
                    int_mem_i [8'hb5] <=  8'hd5 ;
                    int_mem_i [8'hb6] <=  8'h4e ;
                    int_mem_i [8'hb7] <=  8'ha9 ;
                    int_mem_i [8'hb8] <=  8'h6c ;
                    int_mem_i [8'hb9] <=  8'h56 ;
                    int_mem_i [8'hba] <=  8'hf4 ;
                    int_mem_i [8'hbb] <=  8'hea ;
                    int_mem_i [8'hbc] <=  8'h65 ;
                    int_mem_i [8'hbd] <=  8'h7a ;
                    int_mem_i [8'hbe] <=  8'hae ;
                    int_mem_i [8'hbf] <=  8'h08 ;
                    int_mem_i [8'hc0] <=  8'hba ;
                    int_mem_i [8'hc1] <=  8'h78 ;
                    int_mem_i [8'hc2] <=  8'h25 ;
                    int_mem_i [8'hc3] <=  8'h2e ;
                    int_mem_i [8'hc4] <=  8'h1c ;
                    int_mem_i [8'hc5] <=  8'ha6 ;
                    int_mem_i [8'hc6] <=  8'hb4 ;
                    int_mem_i [8'hc7] <=  8'hc6 ;
                    int_mem_i [8'hc8] <=  8'he8 ;
                    int_mem_i [8'hc9] <=  8'hdd ;
                    int_mem_i [8'hca] <=  8'h74 ;
                    int_mem_i [8'hcb] <=  8'h1f ;
                    int_mem_i [8'hcc] <=  8'h4b ;
                    int_mem_i [8'hcd] <=  8'hbd ;
                    int_mem_i [8'hce] <=  8'h8b ;
                    int_mem_i [8'hcf] <=  8'h8a ;
                    int_mem_i [8'hd0] <=  8'h70 ;
                    int_mem_i [8'hd1] <=  8'h3e ;
                    int_mem_i [8'hd2] <=  8'hb5 ;
                    int_mem_i [8'hd3] <=  8'h66 ;
                    int_mem_i [8'hd4] <=  8'h48 ;
                    int_mem_i [8'hd5] <=  8'h03 ;
                    int_mem_i [8'hd6] <=  8'hf6 ;
                    int_mem_i [8'hd7] <=  8'h0e ;
                    int_mem_i [8'hd8] <=  8'h61 ;
                    int_mem_i [8'hd9] <=  8'h35 ;
                    int_mem_i [8'hda] <=  8'h57 ;
                    int_mem_i [8'hdb] <=  8'hb9 ;
                    int_mem_i [8'hdc] <=  8'h86 ;
                    int_mem_i [8'hdd] <=  8'hc1 ;
                    int_mem_i [8'hde] <=  8'h1d ;
                    int_mem_i [8'hdf] <=  8'h9e ;
                    int_mem_i [8'he0] <=  8'he1 ;
                    int_mem_i [8'he1] <=  8'hf8 ;
                    int_mem_i [8'he2] <=  8'h98 ;
                    int_mem_i [8'he3] <=  8'h11 ;
                    int_mem_i [8'he4] <=  8'h69 ;
                    int_mem_i [8'he5] <=  8'hd9 ;
                    int_mem_i [8'he6] <=  8'h8e ;
                    int_mem_i [8'he7] <=  8'h94 ;
                    int_mem_i [8'he8] <=  8'h9b ;
                    int_mem_i [8'he9] <=  8'h1e ;
                    int_mem_i [8'hea] <=  8'h87 ;
                    int_mem_i [8'heb] <=  8'he9 ;
                    int_mem_i [8'hec] <=  8'hce ;
                    int_mem_i [8'hed] <=  8'h55 ;
                    int_mem_i [8'hee] <=  8'h28 ;
                    int_mem_i [8'hef] <=  8'hdf ;
                    int_mem_i [8'hf0] <=  8'h8c ;
                    int_mem_i [8'hf1] <=  8'ha1 ;
                    int_mem_i [8'hf2] <=  8'h89 ;
                    int_mem_i [8'hf3] <=  8'h0d ;
                    int_mem_i [8'hf4] <=  8'hbf ;
                    int_mem_i [8'hf5] <=  8'he6 ;
                    int_mem_i [8'hf6] <=  8'h42 ;
                    int_mem_i [8'hf7] <=  8'h68 ;
                    int_mem_i [8'hf8] <=  8'h41 ;
                    int_mem_i [8'hf9] <=  8'h99 ;
                    int_mem_i [8'hfa] <=  8'h2d ;
                    int_mem_i [8'hfb] <=  8'h0f ;
                    int_mem_i [8'hfc] <=  8'hb0 ;
                    int_mem_i [8'hfd] <=  8'h54 ;
                    int_mem_i [8'hfe] <=  8'hbb ;
                    int_mem_i [8'hff] <=  8'h16 ;
        end
		else begin
			mem_out= int_mem_i[ad];
		end
	end
endmodule 



